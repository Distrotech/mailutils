if address :is :all "from" "tim@example.com" {
  discard;
}

