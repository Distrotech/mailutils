if header :contains ["from"] ["idiot@example.edu"]
  {
    discard;
  }
