if exists "X"
  {
    keep;
  }

