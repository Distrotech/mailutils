if size :over 100K { /* this is a comment
  this is still a comment */ discard /* this is a comment
    */ ;
}
