# -*- sieve -*-
# This file is part of Mailutils testsuite.
# Copyright (C) 2002, Free Software Foundation.
# See file COPYING for distribution conditions.

if header ["X-Caffeine","Subject"] ["C8H10N4O2","Coffee"] {
        discard;
}

