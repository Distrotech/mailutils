if size :under 1M { keep; } else { discard; }

