require "fileinto";

if exists "subject"
{
    fileinto "subject";
}

