
  if not size :under 1M { discard; }

