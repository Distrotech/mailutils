# an empty script

