require ["fileinto", "reject"];
require "fileinto";
# require "vacation";

