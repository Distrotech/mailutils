# -*- sieve -*-
# This file is part of Mailutils testsuite.
# Copyright (C) 2002, 2007 Free Software Foundation.
# See file COPYING for distribution conditions.

require "fileinto";

fileinto "+file";
