if exists "X"
{
    keep;
}

