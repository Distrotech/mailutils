
require "fileinto";

fileinto "./_save-all.mbox";

