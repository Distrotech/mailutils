if size :under 500K {
    discard;
}

keep;
