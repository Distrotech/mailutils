  if header :contains :comparator "i;octet" "Subject"
                "MAKE MONEY FAST" {
                   discard;
             }

