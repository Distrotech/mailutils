  if size :over 550 { # this is a comment
      discard;
  }
