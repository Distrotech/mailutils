require "envelope";

if envelope :all :is "from" "tim@example.com"
  {
    discard;
  }
