# -*- sieve -*-
# This file is part of Mailutils testsuite.
# Copyright (C) 2002, Free Software Foundation.
# See file COPYING for distribution conditions.

require "fileinto";

if address :localpart :is ["To", "Cc"] [ "foo", "oof" ]
  {
    discard;
  } 
